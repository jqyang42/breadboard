module register_65(outA, clk, ie, oeA, clr, in, write_ctrl);
    input clk, ie, oeA, clr, write_ctrl;
    input [64:0] in;

    output [64:0] outA;
    
    wire [64:0] dff_out;

    and input_enable(w_ie, ie, write_ctrl);

    dffe_ref dffe0(.q(dff_out[0]), .d(in[0]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe1(.q(dff_out[1]), .d(in[1]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe2(.q(dff_out[2]), .d(in[2]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe3(.q(dff_out[3]), .d(in[3]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe4(.q(dff_out[4]), .d(in[4]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe5(.q(dff_out[5]), .d(in[5]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe6(.q(dff_out[6]), .d(in[6]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe7(.q(dff_out[7]), .d(in[7]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe8(.q(dff_out[8]), .d(in[8]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe9(.q(dff_out[9]), .d(in[9]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe10(.q(dff_out[10]), .d(in[10]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe11(.q(dff_out[11]), .d(in[11]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe12(.q(dff_out[12]), .d(in[12]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe13(.q(dff_out[13]), .d(in[13]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe14(.q(dff_out[14]), .d(in[14]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe15(.q(dff_out[15]), .d(in[15]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe16(.q(dff_out[16]), .d(in[16]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe17(.q(dff_out[17]), .d(in[17]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe18(.q(dff_out[18]), .d(in[18]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe19(.q(dff_out[19]), .d(in[19]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe20(.q(dff_out[20]), .d(in[20]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe21(.q(dff_out[21]), .d(in[21]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe22(.q(dff_out[22]), .d(in[22]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe23(.q(dff_out[23]), .d(in[23]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe24(.q(dff_out[24]), .d(in[24]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe25(.q(dff_out[25]), .d(in[25]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe26(.q(dff_out[26]), .d(in[26]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe27(.q(dff_out[27]), .d(in[27]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe28(.q(dff_out[28]), .d(in[28]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe29(.q(dff_out[29]), .d(in[29]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe30(.q(dff_out[30]), .d(in[30]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe31(.q(dff_out[31]), .d(in[31]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe32(.q(dff_out[32]), .d(in[32]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe33(.q(dff_out[33]), .d(in[33]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe34(.q(dff_out[34]), .d(in[34]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe35(.q(dff_out[35]), .d(in[35]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe36(.q(dff_out[36]), .d(in[36]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe37(.q(dff_out[37]), .d(in[37]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe38(.q(dff_out[38]), .d(in[38]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe39(.q(dff_out[39]), .d(in[39]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe40(.q(dff_out[40]), .d(in[40]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe41(.q(dff_out[41]), .d(in[41]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe42(.q(dff_out[42]), .d(in[42]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe43(.q(dff_out[43]), .d(in[43]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe44(.q(dff_out[44]), .d(in[44]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe45(.q(dff_out[45]), .d(in[45]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe46(.q(dff_out[46]), .d(in[46]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe47(.q(dff_out[47]), .d(in[47]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe48(.q(dff_out[48]), .d(in[48]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe49(.q(dff_out[49]), .d(in[49]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe50(.q(dff_out[50]), .d(in[50]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe51(.q(dff_out[51]), .d(in[51]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe52(.q(dff_out[52]), .d(in[52]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe53(.q(dff_out[53]), .d(in[53]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe54(.q(dff_out[54]), .d(in[54]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe55(.q(dff_out[55]), .d(in[55]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe56(.q(dff_out[56]), .d(in[56]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe57(.q(dff_out[57]), .d(in[57]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe58(.q(dff_out[58]), .d(in[58]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe59(.q(dff_out[59]), .d(in[59]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe60(.q(dff_out[60]), .d(in[60]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe61(.q(dff_out[61]), .d(in[61]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe62(.q(dff_out[62]), .d(in[62]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe63(.q(dff_out[63]), .d(in[63]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe64(.q(dff_out[64]), .d(in[64]), .clk(clk), .en(w_ie), .clr(clr));

    tri_state outputA0(.out(outA[0]), .in(dff_out[0]), .oe(oeA));
    tri_state outputA1(.out(outA[1]), .in(dff_out[1]), .oe(oeA));
    tri_state outputA2(.out(outA[2]), .in(dff_out[2]), .oe(oeA));
    tri_state outputA3(.out(outA[3]), .in(dff_out[3]), .oe(oeA));
    tri_state outputA4(.out(outA[4]), .in(dff_out[4]), .oe(oeA));
    tri_state outputA5(.out(outA[5]), .in(dff_out[5]), .oe(oeA));
    tri_state outputA6(.out(outA[6]), .in(dff_out[6]), .oe(oeA));
    tri_state outputA7(.out(outA[7]), .in(dff_out[7]), .oe(oeA));
    tri_state outputA8(.out(outA[8]), .in(dff_out[8]), .oe(oeA));
    tri_state outputA9(.out(outA[9]), .in(dff_out[9]), .oe(oeA));
    tri_state outputA10(.out(outA[10]), .in(dff_out[10]), .oe(oeA));
    tri_state outputA11(.out(outA[11]), .in(dff_out[11]), .oe(oeA));
    tri_state outputA12(.out(outA[12]), .in(dff_out[12]), .oe(oeA));
    tri_state outputA13(.out(outA[13]), .in(dff_out[13]), .oe(oeA));
    tri_state outputA14(.out(outA[14]), .in(dff_out[14]), .oe(oeA));
    tri_state outputA15(.out(outA[15]), .in(dff_out[15]), .oe(oeA));
    tri_state outputA16(.out(outA[16]), .in(dff_out[16]), .oe(oeA));
    tri_state outputA17(.out(outA[17]), .in(dff_out[17]), .oe(oeA));
    tri_state outputA18(.out(outA[18]), .in(dff_out[18]), .oe(oeA));
    tri_state outputA19(.out(outA[19]), .in(dff_out[19]), .oe(oeA));
    tri_state outputA20(.out(outA[20]), .in(dff_out[20]), .oe(oeA));
    tri_state outputA21(.out(outA[21]), .in(dff_out[21]), .oe(oeA));
    tri_state outputA22(.out(outA[22]), .in(dff_out[22]), .oe(oeA));
    tri_state outputA23(.out(outA[23]), .in(dff_out[23]), .oe(oeA));
    tri_state outputA24(.out(outA[24]), .in(dff_out[24]), .oe(oeA));
    tri_state outputA25(.out(outA[25]), .in(dff_out[25]), .oe(oeA));
    tri_state outputA26(.out(outA[26]), .in(dff_out[26]), .oe(oeA));
    tri_state outputA27(.out(outA[27]), .in(dff_out[27]), .oe(oeA));
    tri_state outputA28(.out(outA[28]), .in(dff_out[28]), .oe(oeA));
    tri_state outputA29(.out(outA[29]), .in(dff_out[29]), .oe(oeA));
    tri_state outputA30(.out(outA[30]), .in(dff_out[30]), .oe(oeA));
    tri_state outputA31(.out(outA[31]), .in(dff_out[31]), .oe(oeA));
    tri_state outputA32(.out(outA[32]), .in(dff_out[32]), .oe(oeA));
    tri_state outputA33(.out(outA[33]), .in(dff_out[33]), .oe(oeA));
    tri_state outputA34(.out(outA[34]), .in(dff_out[34]), .oe(oeA));
    tri_state outputA35(.out(outA[35]), .in(dff_out[35]), .oe(oeA));
    tri_state outputA36(.out(outA[36]), .in(dff_out[36]), .oe(oeA));
    tri_state outputA37(.out(outA[37]), .in(dff_out[37]), .oe(oeA));
    tri_state outputA38(.out(outA[38]), .in(dff_out[38]), .oe(oeA));
    tri_state outputA39(.out(outA[39]), .in(dff_out[39]), .oe(oeA));
    tri_state outputA40(.out(outA[40]), .in(dff_out[40]), .oe(oeA));
    tri_state outputA41(.out(outA[41]), .in(dff_out[41]), .oe(oeA));
    tri_state outputA42(.out(outA[42]), .in(dff_out[42]), .oe(oeA));
    tri_state outputA43(.out(outA[43]), .in(dff_out[43]), .oe(oeA));
    tri_state outputA44(.out(outA[44]), .in(dff_out[44]), .oe(oeA));
    tri_state outputA45(.out(outA[45]), .in(dff_out[45]), .oe(oeA));
    tri_state outputA46(.out(outA[46]), .in(dff_out[46]), .oe(oeA));
    tri_state outputA47(.out(outA[47]), .in(dff_out[47]), .oe(oeA));
    tri_state outputA48(.out(outA[48]), .in(dff_out[48]), .oe(oeA));
    tri_state outputA49(.out(outA[49]), .in(dff_out[49]), .oe(oeA));
    tri_state outputA50(.out(outA[50]), .in(dff_out[50]), .oe(oeA));
    tri_state outputA51(.out(outA[51]), .in(dff_out[51]), .oe(oeA));
    tri_state outputA52(.out(outA[52]), .in(dff_out[52]), .oe(oeA));
    tri_state outputA53(.out(outA[53]), .in(dff_out[53]), .oe(oeA));
    tri_state outputA54(.out(outA[54]), .in(dff_out[54]), .oe(oeA));
    tri_state outputA55(.out(outA[55]), .in(dff_out[55]), .oe(oeA));
    tri_state outputA56(.out(outA[56]), .in(dff_out[56]), .oe(oeA));
    tri_state outputA57(.out(outA[57]), .in(dff_out[57]), .oe(oeA));
    tri_state outputA58(.out(outA[58]), .in(dff_out[58]), .oe(oeA));
    tri_state outputA59(.out(outA[59]), .in(dff_out[59]), .oe(oeA));
    tri_state outputA60(.out(outA[60]), .in(dff_out[60]), .oe(oeA));
    tri_state outputA61(.out(outA[61]), .in(dff_out[61]), .oe(oeA));
    tri_state outputA62(.out(outA[62]), .in(dff_out[62]), .oe(oeA));
    tri_state outputA63(.out(outA[63]), .in(dff_out[63]), .oe(oeA));
    tri_state outputA64(.out(outA[64]), .in(dff_out[64]), .oe(oeA));
endmodule