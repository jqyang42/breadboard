module or_gate(A, B, out);
    input [31:0] A, B;
    output [31:0] out;

    or gate0(out[0], A[0], B[0]);
    or gate1(out[1], A[1], B[1]);
    or gate2(out[2], A[2], B[2]);
    or gate3(out[3], A[3], B[3]);
    or gate4(out[4], A[4], B[4]);
    or gate5(out[5], A[5], B[5]);
    or gate6(out[6], A[6], B[6]);
    or gate7(out[7], A[7], B[7]);
    or gate8(out[8], A[8], B[8]);
    or gate9(out[9], A[9], B[9]);
    or gate10(out[10], A[10], B[10]);
    or gate11(out[11], A[11], B[11]);
    or gate12(out[12], A[12], B[12]);
    or gate13(out[13], A[13], B[13]);
    or gate14(out[14], A[14], B[14]);
    or gate15(out[15], A[15], B[15]);
    or gate16(out[16], A[16], B[16]);
    or gate17(out[17], A[17], B[17]);
    or gate18(out[18], A[18], B[18]);
    or gate19(out[19], A[19], B[19]);
    or gate20(out[20], A[20], B[20]);
    or gate21(out[21], A[21], B[21]);
    or gate22(out[22], A[22], B[22]);
    or gate23(out[23], A[23], B[23]);
    or gate24(out[24], A[24], B[24]);
    or gate25(out[25], A[25], B[25]);
    or gate26(out[26], A[26], B[26]);
    or gate27(out[27], A[27], B[27]);
    or gate28(out[28], A[28], B[28]);
    or gate29(out[29], A[29], B[29]);
    or gate30(out[30], A[30], B[30]);
    or gate31(out[31], A[31], B[31]);
endmodule