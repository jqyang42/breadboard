module register_32(outA, outB, clk, ie, oeA, oeB, clr, in, write_ctrl);
    input clk, ie, oeA, oeB, clr, write_ctrl;
    input [31:0] in;

    output [31:0] outA, outB;
    
    wire [31:0] dff_out;

    and input_enable(w_ie, ie, write_ctrl);

    dffe_ref dffe0(.q(dff_out[0]), .d(in[0]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe1(.q(dff_out[1]), .d(in[1]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe2(.q(dff_out[2]), .d(in[2]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe3(.q(dff_out[3]), .d(in[3]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe4(.q(dff_out[4]), .d(in[4]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe5(.q(dff_out[5]), .d(in[5]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe6(.q(dff_out[6]), .d(in[6]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe7(.q(dff_out[7]), .d(in[7]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe8(.q(dff_out[8]), .d(in[8]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe9(.q(dff_out[9]), .d(in[9]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe10(.q(dff_out[10]), .d(in[10]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe11(.q(dff_out[11]), .d(in[11]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe12(.q(dff_out[12]), .d(in[12]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe13(.q(dff_out[13]), .d(in[13]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe14(.q(dff_out[14]), .d(in[14]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe15(.q(dff_out[15]), .d(in[15]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe16(.q(dff_out[16]), .d(in[16]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe17(.q(dff_out[17]), .d(in[17]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe18(.q(dff_out[18]), .d(in[18]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe19(.q(dff_out[19]), .d(in[19]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe20(.q(dff_out[20]), .d(in[20]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe21(.q(dff_out[21]), .d(in[21]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe22(.q(dff_out[22]), .d(in[22]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe23(.q(dff_out[23]), .d(in[23]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe24(.q(dff_out[24]), .d(in[24]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe25(.q(dff_out[25]), .d(in[25]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe26(.q(dff_out[26]), .d(in[26]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe27(.q(dff_out[27]), .d(in[27]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe28(.q(dff_out[28]), .d(in[28]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe29(.q(dff_out[29]), .d(in[29]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe30(.q(dff_out[30]), .d(in[30]), .clk(clk), .en(w_ie), .clr(clr));
    dffe_ref dffe31(.q(dff_out[31]), .d(in[31]), .clk(clk), .en(w_ie), .clr(clr));

    tri_state outputA0(.out(outA[0]), .in(dff_out[0]), .oe(oeA));
    tri_state outputA1(.out(outA[1]), .in(dff_out[1]), .oe(oeA));
    tri_state outputA2(.out(outA[2]), .in(dff_out[2]), .oe(oeA));
    tri_state outputA3(.out(outA[3]), .in(dff_out[3]), .oe(oeA));
    tri_state outputA4(.out(outA[4]), .in(dff_out[4]), .oe(oeA));
    tri_state outputA5(.out(outA[5]), .in(dff_out[5]), .oe(oeA));
    tri_state outputA6(.out(outA[6]), .in(dff_out[6]), .oe(oeA));
    tri_state outputA7(.out(outA[7]), .in(dff_out[7]), .oe(oeA));
    tri_state outputA8(.out(outA[8]), .in(dff_out[8]), .oe(oeA));
    tri_state outputA9(.out(outA[9]), .in(dff_out[9]), .oe(oeA));
    tri_state outputA10(.out(outA[10]), .in(dff_out[10]), .oe(oeA));
    tri_state outputA11(.out(outA[11]), .in(dff_out[11]), .oe(oeA));
    tri_state outputA12(.out(outA[12]), .in(dff_out[12]), .oe(oeA));
    tri_state outputA13(.out(outA[13]), .in(dff_out[13]), .oe(oeA));
    tri_state outputA14(.out(outA[14]), .in(dff_out[14]), .oe(oeA));
    tri_state outputA15(.out(outA[15]), .in(dff_out[15]), .oe(oeA));
    tri_state outputA16(.out(outA[16]), .in(dff_out[16]), .oe(oeA));
    tri_state outputA17(.out(outA[17]), .in(dff_out[17]), .oe(oeA));
    tri_state outputA18(.out(outA[18]), .in(dff_out[18]), .oe(oeA));
    tri_state outputA19(.out(outA[19]), .in(dff_out[19]), .oe(oeA));
    tri_state outputA20(.out(outA[20]), .in(dff_out[20]), .oe(oeA));
    tri_state outputA21(.out(outA[21]), .in(dff_out[21]), .oe(oeA));
    tri_state outputA22(.out(outA[22]), .in(dff_out[22]), .oe(oeA));
    tri_state outputA23(.out(outA[23]), .in(dff_out[23]), .oe(oeA));
    tri_state outputA24(.out(outA[24]), .in(dff_out[24]), .oe(oeA));
    tri_state outputA25(.out(outA[25]), .in(dff_out[25]), .oe(oeA));
    tri_state outputA26(.out(outA[26]), .in(dff_out[26]), .oe(oeA));
    tri_state outputA27(.out(outA[27]), .in(dff_out[27]), .oe(oeA));
    tri_state outputA28(.out(outA[28]), .in(dff_out[28]), .oe(oeA));
    tri_state outputA29(.out(outA[29]), .in(dff_out[29]), .oe(oeA));
    tri_state outputA30(.out(outA[30]), .in(dff_out[30]), .oe(oeA));
    tri_state outputA31(.out(outA[31]), .in(dff_out[31]), .oe(oeA));

    tri_state outputB0(.out(outB[0]), .in(dff_out[0]), .oe(oeB));
    tri_state outputB1(.out(outB[1]), .in(dff_out[1]), .oe(oeB));
    tri_state outputB2(.out(outB[2]), .in(dff_out[2]), .oe(oeB));
    tri_state outputB3(.out(outB[3]), .in(dff_out[3]), .oe(oeB));
    tri_state outputB4(.out(outB[4]), .in(dff_out[4]), .oe(oeB));
    tri_state outputB5(.out(outB[5]), .in(dff_out[5]), .oe(oeB));
    tri_state outputB6(.out(outB[6]), .in(dff_out[6]), .oe(oeB));
    tri_state outputB7(.out(outB[7]), .in(dff_out[7]), .oe(oeB));
    tri_state outputB8(.out(outB[8]), .in(dff_out[8]), .oe(oeB));
    tri_state outputB9(.out(outB[9]), .in(dff_out[9]), .oe(oeB));
    tri_state outputB10(.out(outB[10]), .in(dff_out[10]), .oe(oeB));
    tri_state outputB11(.out(outB[11]), .in(dff_out[11]), .oe(oeB));
    tri_state outputB12(.out(outB[12]), .in(dff_out[12]), .oe(oeB));
    tri_state outputB13(.out(outB[13]), .in(dff_out[13]), .oe(oeB));
    tri_state outputB14(.out(outB[14]), .in(dff_out[14]), .oe(oeB));
    tri_state outputB15(.out(outB[15]), .in(dff_out[15]), .oe(oeB));
    tri_state outputB16(.out(outB[16]), .in(dff_out[16]), .oe(oeB));
    tri_state outputB17(.out(outB[17]), .in(dff_out[17]), .oe(oeB));
    tri_state outputB18(.out(outB[18]), .in(dff_out[18]), .oe(oeB));
    tri_state outputB19(.out(outB[19]), .in(dff_out[19]), .oe(oeB));
    tri_state outputB20(.out(outB[20]), .in(dff_out[20]), .oe(oeB));
    tri_state outputB21(.out(outB[21]), .in(dff_out[21]), .oe(oeB));
    tri_state outputB22(.out(outB[22]), .in(dff_out[22]), .oe(oeB));
    tri_state outputB23(.out(outB[23]), .in(dff_out[23]), .oe(oeB));
    tri_state outputB24(.out(outB[24]), .in(dff_out[24]), .oe(oeB));
    tri_state outputB25(.out(outB[25]), .in(dff_out[25]), .oe(oeB));
    tri_state outputB26(.out(outB[26]), .in(dff_out[26]), .oe(oeB));
    tri_state outputB27(.out(outB[27]), .in(dff_out[27]), .oe(oeB));
    tri_state outputB28(.out(outB[28]), .in(dff_out[28]), .oe(oeB));
    tri_state outputB29(.out(outB[29]), .in(dff_out[29]), .oe(oeB));
    tri_state outputB30(.out(outB[30]), .in(dff_out[30]), .oe(oeB));
    tri_state outputB31(.out(outB[31]), .in(dff_out[31]), .oe(oeB));
endmodule