module not_gate(A, out);
    input [31:0] A;
    output [31:0] out;

    not not0(out[0], A[0]);
    not not1(out[1], A[1]);
    not not2(out[2], A[2]);
    not not3(out[3], A[3]);
    not not4(out[4], A[4]);
    not not5(out[5], A[5]);
    not not6(out[6], A[6]);
    not not7(out[7], A[7]);
    not not8(out[8], A[8]);
    not not9(out[9], A[9]);
    not not10(out[10], A[10]);
    not not11(out[11], A[11]);
    not not12(out[12], A[12]);
    not not13(out[13], A[13]);
    not not14(out[14], A[14]);
    not not15(out[15], A[15]);
    not not16(out[16], A[16]);
    not not17(out[17], A[17]);
    not not18(out[18], A[18]);
    not not19(out[19], A[19]);
    not not20(out[20], A[20]);
    not not21(out[21], A[21]);
    not not22(out[22], A[22]);
    not not23(out[23], A[23]);
    not not24(out[24], A[24]);
    not not25(out[25], A[25]);
    not not26(out[26], A[26]);
    not not27(out[27], A[27]);
    not not28(out[28], A[28]);
    not not29(out[29], A[29]);
    not not30(out[30], A[30]);
    not not31(out[31], A[31]);
endmodule